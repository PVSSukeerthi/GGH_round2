module rtl1(input A, B, output Y);
    assign Y = A & B;
endmodule

