module rtl8 (input [1:0] A, B, output [3:0] P);
    assign P = A * B;
endmodule

